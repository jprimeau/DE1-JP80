library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;
    
use work.jp80_pkg.all;
    
entity JP80_FILEREG is
    port (
        clk             : in t_wire;
        data_in_h       : in t_data;
        data_in_l       : in t_data;
        we_h            : in t_wire;
        we_l            : in t_wire;
        reg_addr_in     : in t_regaddr;
        reg_addr_out_a  : in t_regaddr;
        reg_addr_out_b  : in t_regaddr;
        data_out_a_h    : out t_data;
        data_out_a_l    : out t_data;
        en_a_h          : in t_wire;
        en_a_l          : in t_wire;
        data_out_b_h    : out t_data;
        data_out_b_l    : out t_data;
        en_b_h          : in t_wire;
        en_b_l          : in t_wire
    );
end JP80_FILEREG;

architecture rtl of JP80_FILEREG is
    type file_register is array(0 to 3) of t_data;
    signal regs_h : file_register;
    signal regs_l : file_register;
begin
    process (clk)
    begin
        if clk'event and clk = '0' then
            if we_h = '1' then
                regs_h(conv_integer(reg_addr_in)) <= data_in_h;
            end if;
            if we_l = '1' then
                regs_l(conv_integer(reg_addr_in)) <= data_in_l;
            end if;
        end if;
    end process;
    data_out_a_h <= regs_h(conv_integer(reg_addr_out_a)) when en_a_h = '1' else (others=>'Z');
    data_out_a_l <= regs_l(conv_integer(reg_addr_out_a)) when en_a_l = '1' else (others=>'Z');
    data_out_b_h <= regs_h(conv_integer(reg_addr_out_b)) when en_b_h = '1' else (others=>'Z');
    data_out_b_l <= regs_l(conv_integer(reg_addr_out_b)) when en_b_l = '1' else (others=>'Z');
end architecture;